LIBRARY ieee;
USE ieee.std_logic_1164.all; 

package constants is

constant NUM_OF_PWMMOD  : natural :=3;

end package constants;
