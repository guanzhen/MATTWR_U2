MAX_OSC_inst : MAX_OSC PORT MAP (
		oscena	 => oscena_sig,
		osc	 => osc_sig
	);
