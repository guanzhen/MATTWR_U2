-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.1.0 Build 162 10/23/2013 SJ Full Version"
-- CREATED		"Fri Oct 13 09:51:24 2017"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY MaterialTowerCPLD IS 
	PORT
	(
		nRD :  IN  STD_LOGIC;
		nWR :  IN  STD_LOGIC;
		nCS :  IN  STD_LOGIC;
		nADV :  IN  STD_LOGIC;
		nWAIT :  IN  STD_LOGIC;
		ENC_1_A :  IN  STD_LOGIC;
		Clk :  IN  STD_LOGIC;
		ENC_1_B :  IN  STD_LOGIC;
		ENC_1_N :  IN  STD_LOGIC;
		ENC_2_A :  IN  STD_LOGIC;
		ENC_2_B :  IN  STD_LOGIC;
		ENC_2_N :  IN  STD_LOGIC;
		PWM_LED :  IN  STD_LOGIC;
		CC_CAN1_TXD :  IN  STD_LOGIC;
		CC_CAN2_TXD :  IN  STD_LOGIC;
		CAN1_RXD :  IN  STD_LOGIC;
		CAN2_RXD :  IN  STD_LOGIC;
		EN_EDIF_CAN :  IN  STD_LOGIC;
		FAN_PULSE :  IN  STD_LOGIC;
		SDCLKO :  IN  STD_LOGIC;
		CPLD_INT :  IN  STD_LOGIC;
		RST :  IN  STD_LOGIC;
		A :  IN  STD_LOGIC_VECTOR(6 DOWNTO 0);
		AD :  INOUT  STD_LOGIC_VECTOR(7 DOWNTO 0);
		DIP_SWITCH :  IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		IO_Input13 :  IN  STD_LOGIC;
		IO_Input12 :  IN  STD_LOGIC;
		IO_Input11 :  IN  STD_LOGIC;
		IO_Input10 :  IN  STD_LOGIC;
		IO_Input9 :  IN  STD_LOGIC;
		IO_Input8 :  IN  STD_LOGIC;
		IO_Input23 :  IN  STD_LOGIC;
		IO_Input22 :  IN  STD_LOGIC;
		IO_Input21 :  IN  STD_LOGIC;
		IO_Input20 :  IN  STD_LOGIC;
		IO_Input19 :  IN  STD_LOGIC;
		IO_Input18 :  IN  STD_LOGIC;
		IO_Input17 :  IN  STD_LOGIC;
		IO_Input16 :  IN  STD_LOGIC;
		IO_Input2 :  IN  STD_LOGIC;
		IO_Input1 :  IN  STD_LOGIC;
		IO_Input0 :  IN  STD_LOGIC;
		ENC_1_PS :  OUT  STD_LOGIC;
		ENC_1_DIR :  OUT  STD_LOGIC;
		ENC_1_INX :  OUT  STD_LOGIC;
		ENC_2_PS :  OUT  STD_LOGIC;
		ENC_2_DIR :  OUT  STD_LOGIC;
		ENC_2_INX :  OUT  STD_LOGIC;
		CAN1_TXD :  OUT  STD_LOGIC;
		CAN2_TXD :  OUT  STD_LOGIC;
		CC_CAN1_RXD :  OUT  STD_LOGIC;
		CC_CAN2_RXD :  OUT  STD_LOGIC;
		ENC_ERR :  OUT  STD_LOGIC;
		FPGA_OK :  OUT  STD_LOGIC;
		FAN_PWM :  OUT  STD_LOGIC;
		LED_PWM :  OUT  STD_LOGIC;
		PIZZA_CALIBRATION :  OUT  STD_LOGIC;
		IO_Output :  OUT  STD_LOGIC_VECTOR(16 DOWNTO 0);
		Seg_LED :  OUT  STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END MaterialTowerCPLD;

ARCHITECTURE bdf_type OF MaterialTowerCPLD IS 

COMPONENT sram_io
GENERIC (CPLD_VERSION : STD_LOGIC_VECTOR(7 DOWNTO 0);
			WIDTH : INTEGER
			);
	PORT(nRESET : IN STD_LOGIC;
		 nRD : IN STD_LOGIC;
		 nWR : IN STD_LOGIC;
		 nCS : IN STD_LOGIC;
		 nADV : IN STD_LOGIC;
		 nWAIT : IN STD_LOGIC;
		 DATA : INOUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 IO_DATA : INOUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 IO_RDY_WR : OUT STD_LOGIC;
		 IO_RDY_RD : OUT STD_LOGIC;
		 IO_RDY_ADR : OUT STD_LOGIC;
		 IO_ADDR : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT io_space
GENERIC (BUS_WIDTH : INTEGER;
			CPLD_VERSION : STD_LOGIC_VECTOR(7 DOWNTO 0);
			ENC_WIDTH : INTEGER;
			FAN_WIDTH : INTEGER
			);
	PORT(nRESET : IN STD_LOGIC;
		 Clk : IN STD_LOGIC;
		 IO_RDY_WR : IN STD_LOGIC;
		 IO_RDY_RD : IN STD_LOGIC;
		 IO_RDY_ADR : IN STD_LOGIC;
		 Seg_DP : IN STD_LOGIC;
		 DIP_SW : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 Enc_MT1 : IN STD_LOGIC_VECTOR(23 DOWNTO 0);
		 Enc_MT2 : IN STD_LOGIC_VECTOR(23 DOWNTO 0);
		 IO_ADDR : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 IO_DATA : INOUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 iPin0_7 : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 iPin16_23 : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 iPin8_15 : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 oPin16_23 : OUT STD_LOGIC;
		 Wr_MT1 : OUT STD_LOGIC;
		 Wr_MT2 : OUT STD_LOGIC;
		 Pizza_Cali : OUT STD_LOGIC;
		 oPin0_7 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 oPin8_15 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 Seg_LED : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
		 WrVal_MT1 : OUT STD_LOGIC_VECTOR(23 DOWNTO 0);
		 WrVal_MT2 : OUT STD_LOGIC_VECTOR(23 DOWNTO 0)
	);
END COMPONENT;

COMPONENT quaddectodirpulse
GENERIC (CPLD_VERSION : STD_LOGIC_VECTOR(7 DOWNTO 0);
			ENC_WIDTH : INTEGER
			);
	PORT(A : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 N : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 Wr : IN STD_LOGIC;
		 WrVal : IN STD_LOGIC_VECTOR(23 DOWNTO 0);
		 PS : OUT STD_LOGIC;
		 DIR : OUT STD_LOGIC;
		 INX : OUT STD_LOGIC;
		 Enc : OUT STD_LOGIC_VECTOR(23 DOWNTO 0)
	);
END COMPONENT;

COMPONENT hex7seg
	PORT(A : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 LED7S : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

SIGNAL	gdfx_temp0 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC_VECTOR(23 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC_VECTOR(23 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC_VECTOR(23 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC_VECTOR(23 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC_VECTOR(4 DOWNTO 0);

SIGNAL	GDFX_TEMP_SIGNAL_0 :  STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_1 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_2 :  STD_LOGIC_VECTOR(5 DOWNTO 0);

BEGIN 
CAN1_TXD <= CC_CAN1_TXD;
CAN2_TXD <= CC_CAN2_TXD;
CC_CAN2_RXD <= CAN2_RXD;
FAN_PWM <= PWM_LED;
LED_PWM <= PWM_LED;
ENC_ERR <= SYNTHESIZED_WIRE_13;

GDFX_TEMP_SIGNAL_0 <= (IO_Input2 & IO_Input1 & IO_Input0);
GDFX_TEMP_SIGNAL_1 <= (IO_Input23 & IO_Input22 & IO_Input21 & IO_Input20 & IO_Input19 & IO_Input18 & IO_Input17 & IO_Input16);
GDFX_TEMP_SIGNAL_2 <= (IO_Input13 & IO_Input12 & IO_Input11 & IO_Input10 & IO_Input9 & IO_Input8);


SYNTHESIZED_WIRE_13 <= RST AND CPLD_INT;


b2v_U2 : sram_io
GENERIC MAP(CPLD_VERSION => "00001101",
			WIDTH => 8
			)
PORT MAP(nRESET => SYNTHESIZED_WIRE_13,
		 nRD => nRD,
		 nWR => nWR,
		 nCS => nCS,
		 nADV => nADV,
		 nWAIT => nWAIT,
		 DATA => AD,
		 IO_DATA => gdfx_temp0,
		 IO_RDY_WR => SYNTHESIZED_WIRE_2,
		 IO_RDY_RD => SYNTHESIZED_WIRE_3,
		 IO_RDY_ADR => SYNTHESIZED_WIRE_4,
		 IO_ADDR => SYNTHESIZED_WIRE_7);


b2v_U3 : io_space
GENERIC MAP(BUS_WIDTH => 8,
			CPLD_VERSION => "00001101",
			ENC_WIDTH => 24,
			FAN_WIDTH => 32
			)
PORT MAP(nRESET => SYNTHESIZED_WIRE_13,
		 Clk => Clk,
		 IO_RDY_WR => SYNTHESIZED_WIRE_2,
		 IO_RDY_RD => SYNTHESIZED_WIRE_3,
		 IO_RDY_ADR => SYNTHESIZED_WIRE_4,
		 Seg_DP => PWM_LED,
		 DIP_SW => DIP_SWITCH,
		 Enc_MT1 => SYNTHESIZED_WIRE_5,
		 Enc_MT2 => SYNTHESIZED_WIRE_6,
		 IO_ADDR => SYNTHESIZED_WIRE_7,
		 IO_DATA => gdfx_temp0,
		 iPin0_7 => GDFX_TEMP_SIGNAL_0,
		 iPin16_23 => GDFX_TEMP_SIGNAL_1,
		 iPin8_15 => GDFX_TEMP_SIGNAL_2,
		 oPin16_23 => IO_Output(16),
		 Wr_MT1 => SYNTHESIZED_WIRE_8,
		 Wr_MT2 => SYNTHESIZED_WIRE_10,
		 Pizza_Cali => PIZZA_CALIBRATION,
		 oPin0_7 => IO_Output(7 DOWNTO 0),
		 oPin8_15 => IO_Output(15 DOWNTO 8),
		 Seg_LED => SYNTHESIZED_WIRE_12,
		 WrVal_MT1 => SYNTHESIZED_WIRE_9,
		 WrVal_MT2 => SYNTHESIZED_WIRE_11);


b2v_U4 : quaddectodirpulse
GENERIC MAP(CPLD_VERSION => "00001101",
			ENC_WIDTH => 24
			)
PORT MAP(A => ENC_1_A,
		 B => ENC_1_B,
		 N => ENC_1_N,
		 CLK => Clk,
		 Wr => SYNTHESIZED_WIRE_8,
		 WrVal => SYNTHESIZED_WIRE_9,
		 PS => ENC_1_PS,
		 DIR => ENC_1_DIR,
		 INX => ENC_1_INX,
		 Enc => SYNTHESIZED_WIRE_5);


b2v_U5 : quaddectodirpulse
GENERIC MAP(CPLD_VERSION => "00001101",
			ENC_WIDTH => 24
			)
PORT MAP(A => ENC_2_A,
		 B => ENC_2_B,
		 N => ENC_2_N,
		 CLK => Clk,
		 Wr => SYNTHESIZED_WIRE_10,
		 WrVal => SYNTHESIZED_WIRE_11,
		 PS => ENC_2_PS,
		 DIR => ENC_2_DIR,
		 INX => ENC_2_INX,
		 Enc => SYNTHESIZED_WIRE_6);


b2v_U6 : hex7seg
PORT MAP(A => SYNTHESIZED_WIRE_12,
		 LED7S => Seg_LED);


FPGA_OK <= NOT(Clk AND PWM_LED);


PROCESS(CAN1_RXD,EN_EDIF_CAN)
BEGIN
if (EN_EDIF_CAN = '1') THEN
	CC_CAN1_RXD <= CAN1_RXD;
ELSE
	CC_CAN1_RXD <= 'Z';
END IF;
END PROCESS;


END bdf_type;